* Qucs 0.0.21 /home/saul/projects/QUCS/QUCS_ANALOG_ELEKTRONIK/IE1202_F2_prj/komparator_ngspice.sch
.INCLUDE "/usr/local/share/qucs-s/xspice_cmlib/include/ngspice_mathfunc.inc"
* Qucs 0.0.21  /home/saul/projects/QUCS/QUCS_ANALOG_ELEKTRONIK/IE1202_F2_prj/komparator_ngspice.sch

.SUBCKT Ideal_OpAmp gnd in_p in_m out AOLDC=106 GBP=1e6 RO=75 VLIMP=14 VLIMN=-14 
.PARAM OLG = {10**(AOLDC/20)}
.PARAM Fg = {GBP/OLG}
.PARAM pi = 3.14159
.PARAM C1 = {1e-3/sqrt(2*pi*fg)}
.PARAM R1 = {1e3/sqrt(2*pi*fg)}
ESRC1 _net0 0 in_p in_m OLG
R2 out  _net1 RO
R1 nC  _net0 R1
C1 nC  0 C1
B1 _net1  0  V = V(nC)*u(VLIMP-V(nC))*u(V(nC)-VLIMN)+VLIMP*u(V(nC)-VLIMP)+VLIMN*u(VLIMN-V(nC)) 
.ENDS
           

XOP1 0  Uin Ut Uut Ideal_OpAmp GBP=1E6 AOLDC=106 RO=75 VLIMP=14 VLIMN=-14
V2 Uin 0 DC {V_IN}
V1 Ut 0 DC 5
.control
echo "" > spice4qucs.cir.noise
echo "" > spice4qucs.cir.pz
dc v_in -14 14 0.0996441
write komparator_ngspice_dc.txt v(Uin) v(Ut) v(Uut) 
destroy all
reset

exit
.endc
.END
