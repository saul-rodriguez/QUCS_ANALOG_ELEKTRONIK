* Qucs 0.0.20 /home/saul/projects/QUCS/QUCS_ANALOG_ELEKTRONIK/IE1202_HEMLAB_prj/F11_LAB1_NGSPICE.sch
.INCLUDE "/usr/local/share/qucs-s/xspice_cmlib/include/ngspice_mathfunc.inc"
* Qucs 0.0.20  /home/saul/projects/QUCS/QUCS_ANALOG_ELEKTRONIK/IE1202_HEMLAB_prj/F11_LAB1_NGSPICE.sch
.INCLUDE "/home/saul/projects/QUCS/QUCS_ANALOG_ELEKTRONIK/IE1202_HEMLAB_prj/bcmodels.lib"
.PARAM VIN=1
VPr1 _net0 _net1 DC 0
VPr5 _net2 0 DC 0
VPr4 _net0 _net3 DC 0
R1 B _net3  22000
V1 _net0 0 DC 5
R2 0 B  5600
C2 B _net4  10U 
V3 _net4 0 DC 0 SIN(0 {VIN} 1K 0 0) AC {VIN}
Q1 C  B  E  bc547c

R5 _net2 E  200
R4 C _net1  1000
.control
echo "" > spice4qucs.cir.noise
echo "" > spice4qucs.cir.pz
*let VIN=1
*let VIN=0.01
*ac dec 11 1 10meg 
*write F11_LAB1_NGSPICE_ac.txt v(B) v(C) v(E) VPr1#branch VPr4#branch VPr5#branch 
*destroy all
*reset

*let VIN=1
*let VIN=0.01
*tran 9.999e-08 0.001 0 
*write F11_LAB1_NGSPICE_tran.txt v(B) v(C) v(E) VPr1#branch VPr4#branch VPr5#branch 
*destroy all
*reset
*exit
op
show all

.endc
.END
