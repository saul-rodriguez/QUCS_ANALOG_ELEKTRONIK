* Qucs 0.0.21 /home/saul/projects/QUCS/QUCS_ANALOG_ELEKTRONIK/IE1202_F7_prj/diode_res_tran_ngspice.sch
.INCLUDE "/usr/local/share/qucs-s/xspice_cmlib/include/ngspice_mathfunc.inc"
* Qucs 0.0.21  /home/saul/projects/QUCS/QUCS_ANALOG_ELEKTRONIK/IE1202_F7_prj/diode_res_tran_ngspice.sch
.PARAM V=0.732-0.725
.PARAM I=6.22m-5.34m
.PARAM R=V/I=7.95
VPr1 _net0 Vd DC 0
D_1N4148_1 Vd 0 DMOD_D_1N4148_1 AREA=1.0 Temp=26.85
.MODEL DMOD_D_1N4148_1 D (Is=2.22e-10 N=1.65 Cj0=4e-12 M=0.333 Vj=0.7 Fc=0.5 Rs=0.0686 Tt=5.76e-09 Ikf=0 Kf=0 Af=1 Bv=75 Ibv=1e-06 Xti=3 Eg=1.11 Tcv=0 Trs=0 Ttt1=0 Ttt2=0 Tm1=0 Tm2=0 Tnom=26.85 )
R1 _net1 _net0  220
V1 _net2 0 DC 2
V2 _net1 _net2 DC 0 SIN(0 0.1 1K 0 0 0) AC 0.1
.control
echo "" > spice4qucs.cir.noise
echo "" > spice4qucs.cir.pz
let V=0.732-0.725
let I=6.22m-5.34m
let R=V/I=7.95
tran 9.97506e-06 0.004 0 
write diode_res_tran_ngspice_tran.txt VPr1#branch v(Vd) 
destroy all
reset

exit
.endc
.END
